*** SPICE deck for cell milestone_test{sch} from library Project2
*** Created on Thu Nov 19, 2015 19:37:04
*** Last revised on Sat Nov 21, 2015 17:41:04
*** Written on Sat Nov 21, 2015 18:02:42 by Electric VLSI Design System, 
*version 8.10
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.OPTIONS NOMOD NOPAGE

*** CELL: 6TSRAM{sch}
.SUBCKT _6TSRAM BL BL_B WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@2 WL BL gnd N L=0.022U W=0.22U
Mnmos@1 BL_B WL net@5 gnd N L=0.022U W=0.022U
Mnmos@2 net@5 net@2 gnd gnd N L=0.022U W=0.22U
Mnmos@3 net@2 net@5 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd net@2 net@5 vdd P L=0.022U W=0.22U
Mpmos@1 vdd net@5 net@2 vdd P L=0.022U W=0.022U
.ENDS _6TSRAM

*** CELL: Project1:notBaseline{sch}
.SUBCKT notBaseline in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd in out vdd P L=0.022U W=0.022U
.ENDS notBaseline

*** CELL: precharge{sch}
.SUBCKT precharge BL BL_B Clk_B
** GLOBAL vdd
Mpmos@0 vdd Clk_B BL_B vdd P L=0.022U W=0.022U
Mpmos@1 vdd Clk_B BL vdd P L=0.022U W=0.022U
.ENDS precharge

*** CELL: tri_state_inverter{sch}
.SUBCKT tri_state_inverter En Out data
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@16 En gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@3 data gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@3 En Out gnd N L=0.022U W=0.022U
Mpmos@0 vdd En net@16 vdd P L=0.022U W=0.022U
Mpmos@1 vdd data net@3 vdd P L=0.022U W=0.022U
Mpmos@2 Out net@16 net@3 vdd P L=0.022U W=0.022U
.ENDS tri_state_inverter

*** CELL: milestone{sch}
.SUBCKT milestone Clk_B En Read WL Wdata
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@0 net@88 gnd gnd N L=0.044U W=0.044U
Mpmos@0 vdd net@88 net@0 vdd P L=0.022U W=0.11U
X_6TSRAM@0 net@0 net@4 WL _6TSRAM
XnotBasel@0 En net@46 notBaseline
Xprecharg@0 net@0 net@4 Clk_B precharge
Xtri_stat@2 net@46 Read net@4 tri_state_inverter
Xtri_stat@3 En net@88 Wdata tri_state_inverter
Xtri_stat@5 En net@4 Wdata tri_state_inverter
.ENDS milestone

.global gnd vdd

*** TOP LEVEL CELL: milestone_test{sch}
VVPWL@0 en gnd pwl (0ps 0V 1.5ns 0V 1.6ns 1V 3.2ns 1V 3.3ns 0V 5.5ns 0V 5.6ns 
+1V 7.2ns 1V 7.3ns 0V) DC 0V AC 0V 0
VVPWL@1 wdata gnd pwl (0ps 0V 1.5ns 0V 1.6ns 1V 3.2ns 1V 3.3ns 0V) DC 0V AC 
+0V 0
VVPulse@0 clock gnd pulse (0 1V 0ns 0ps 0ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@1 net@27 gnd pulse (0V 0 0ns 0ps 0ps 1ns 2ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xmileston@0 clock en Read clock wdata milestone
* Trailer cards are described in this file:
.include /home/aasif/Desktop/22nm_HP.pm
.END
