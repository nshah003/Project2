*** SPICE deck for cell size_logic_test{sch} from library Project2
*** Created on Wed Dec 02, 2015 23:12:26
*** Last revised on Thu Dec 03, 2015 03:03:46
*** Written on Thu Dec 03, 2015 03:04:46 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /Users/neilnshah/Desktop/JUNIOR-YEAR/Fall15/Courses/ESE370/Project2/Project2/22nm_HP.pm

*** SUBCIRCUIT Project2__and3 FROM CELL and3{sch}
.SUBCKT Project2__and3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@2 A net@11 gnd N L=0.022U W=0.022U
Mnmos@1 net@11 B net@12 gnd N L=0.022U W=0.022U
Mnmos@2 net@12 C gnd gnd N L=0.022U W=0.022U
Mnmos@3 O net@2 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd C net@2 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@2 O vdd P L=0.022U W=0.022U
Mpmos@2 vdd B net@2 vdd P L=0.022U W=0.022U
Mpmos@3 vdd A net@2 vdd P L=0.022U W=0.022U
.ENDS Project2__and3

*** SUBCIRCUIT Project1__nandBaseline FROM CELL Project1:nandBaseline{sch}
.SUBCKT Project1__nandBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd x out vdd P L=0.022U W=0.022U
Mpmos@1 vdd y out vdd P L=0.022U W=0.022U
.ENDS Project1__nandBaseline

*** SUBCIRCUIT Project1__xorPass FROM CELL Project1:xorPass{sch}
.SUBCKT Project1__xorPass out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@150 y gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@166 net@130 net@150 gnd N L=0.022U W=0.022U
Mnmos@3 y x net@166 gnd N L=0.022U W=0.022U
Mnmos@4 net@130 x gnd gnd N L=0.022U W=0.022U
Mnmos@5 out net@166 gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd y net@150 vdd P L=0.022U W=0.022U
Mpmos@2 vdd x net@130 vdd P L=0.022U W=0.022U
Mpmos@3 vdd net@166 out vdd P L=0.022U W=0.022U
.ENDS Project1__xorPass

*** SUBCIRCUIT Project2__full_adder FROM CELL full_adder{sch}
.SUBCKT Project2__full_adder A B Cin Cout S
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@3 B A Project1__nandBaseline
XnandBase@1 net@16 net@17 Cin Project1__nandBaseline
XnandBase@2 Cout net@3 net@16 Project1__nandBaseline
XxorPass@0 net@17 B A Project1__xorPass
XxorPass@1 S Cin net@17 Project1__xorPass
.ENDS Project2__full_adder

*** SUBCIRCUIT Project2__nor3 FROM CELL nor3{sch}
.SUBCKT Project2__nor3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O C gnd gnd N L=0.022U W=0.022U
Mnmos@1 O B gnd gnd N L=0.022U W=0.022U
Mnmos@2 O A gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A net@0 vdd P L=0.022U W=0.022U
Mpmos@1 net@0 B net@1 vdd P L=0.022U W=0.022U
Mpmos@2 net@1 C O vdd P L=0.022U W=0.022U
.ENDS Project2__nor3

*** SUBCIRCUIT Project1__notBaseline FROM CELL Project1:notBaseline{sch}
.SUBCKT Project1__notBaseline in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd in out vdd P L=0.022U W=0.022U
.ENDS Project1__notBaseline

*** SUBCIRCUIT Project2__size_logic FROM CELL size_logic{sch}
.SUBCKT Project2__size_logic A A_next B B_next C C_next D E Empty Full
** GLOBAL gnd
** GLOBAL vdd
Xand3@0 C_next B_next A_next Full Project2__and3
Xfull_add@0 C net@168 gnd net@158 C_next Project2__full_adder
Xfull_add@1 B net@168 net@158 net@163 B_next Project2__full_adder
Xfull_add@2 A net@187 net@163 full_add@2_Cout A_next Project2__full_adder
XnandBase@0 net@198 D net@199 Project1__nandBaseline
Xnor3@0 C_next B_next A_next Empty Project2__nor3
XnotBasel@3 net@198 net@168 Project1__notBaseline
XnotBasel@4 E net@199 Project1__notBaseline
XxorPass@0 net@187 D E Project1__xorPass
.ENDS Project2__size_logic

.global gnd vdd

*** TOP LEVEL CELL: size_logic_test{sch}
VVPulse@0 D gnd pulse (1V 0V 0ns 0ps 0ps 2ns 4ns) DC 0V AC 0V 0
VVPulse@1 C gnd pulse (1V 0V 0ns 0ps 0ps 4ns 8ns) DC 0V AC 0V 0
VVPulse@2 B gnd pulse (1V 0V 0ns 0ps 0ps 8ns 16ns) DC 0V AC 0V 0
VVPulse@3 A gnd pulse (1V 0V 0ns 0ps 0ps 16ns 32ns) DC 0V AC 0V 0
VVPulse@4 E gnd pulse (1V 0V 0ns 0ps 0ps 1ns 2ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xsize_log@0 A A_next B B_next C C_next D E Empty Full Project2__size_logic
.END
