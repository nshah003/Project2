*** SPICE deck for cell memory_core_test{sch} from library Project2
*** Created on Thu Dec 03, 2015 14:08:13
*** Last revised on Thu Dec 03, 2015 20:18:26
*** Written on Thu Dec 03, 2015 22:19:37 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /Users/neilnshah/Desktop/JUNIOR-YEAR/Fall15/Courses/ESE370/Project2/Project2/22nm_HP.pm

*** SUBCIRCUIT Project1__notBaseline FROM CELL Project1:notBaseline{sch}
.SUBCKT Project1__notBaseline in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd in out vdd P L=0.022U W=0.022U
.ENDS Project1__notBaseline

*** SUBCIRCUIT Project1__nandBaseline FROM CELL Project1:nandBaseline{sch}
.SUBCKT Project1__nandBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd x out vdd P L=0.022U W=0.022U
Mpmos@1 vdd y out vdd P L=0.022U W=0.022U
.ENDS Project1__nandBaseline

*** SUBCIRCUIT HW7__nand_latch FROM CELL HW7:nand_latch{sch}
.SUBCKT HW7__nand_latch clock in out
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@0 in clock Project1__nandBaseline
XnandBase@1 net@11 a out Project1__nandBaseline
XnandBase@2 out net@0 net@11 Project1__nandBaseline
XnotBasel@0 clock a Project1__notBaseline
.ENDS HW7__nand_latch

*** SUBCIRCUIT HW7__register FROM CELL HW7:register{sch}
.SUBCKT HW7__register clock in out
** GLOBAL gnd
** GLOBAL vdd
Xnand_lat@0 clock mid out HW7__nand_latch
Xnand_lat@1 net@17 in mid HW7__nand_latch
XnotBasel@0 clock net@17 Project1__notBaseline
.ENDS HW7__register

*** SUBCIRCUIT Project2__vwide_not FROM CELL vwide_not{sch}
.SUBCKT Project2__vwide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.22U
Mpmos@0 vdd A O vdd P L=0.022U W=0.22U
.ENDS Project2__vwide_not

*** SUBCIRCUIT Project2__clock_div FROM CELL clock_div{sch}
.SUBCKT Project2__clock_div Clk_fast Clk_slow
** GLOBAL gnd
** GLOBAL vdd
XnotBasel@0 net@7 net@4 Project1__notBaseline
Xregister@0 Clk_fast net@4 net@7 HW7__register
Xvwide_no@0 net@4 Clk_slow Project2__vwide_not
.ENDS Project2__clock_div

*** SUBCIRCUIT Project1__norBaseline FROM CELL Project1:norBaseline{sch}
.SUBCKT Project1__norBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x gnd gnd N L=0.022U W=0.022U
Mnmos@1 out y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd y net@10 vdd P L=0.022U W=0.022U
Mpmos@1 net@10 x out vdd P L=0.022U W=0.022U
.ENDS Project1__norBaseline

*** SUBCIRCUIT Project2__wide_not FROM CELL wide_not{sch}
.SUBCKT Project2__wide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.088U
Mpmos@0 vdd A O vdd P L=0.022U W=0.088U
.ENDS Project2__wide_not

*** SUBCIRCUIT Project2__2_4_decoder FROM CELL 2_4_decoder{sch}
.SUBCKT Project2__2_4_decoder B C Clk En WL0 WL1 WL2 WL3
** GLOBAL gnd
** GLOBAL vdd
X_ net@75 net@79 Project1__notBaseline
XnandBase@0 net@73 En net@37 Project1__nandBaseline
XnandBase@1 net@74 En net@36 Project1__nandBaseline
XnandBase@2 net@75 En net@35 Project1__nandBaseline
XnandBase@3 net@76 En net@34 Project1__nandBaseline
XnandBase@4 net@93 Clk net@77 Project1__nandBaseline
XnandBase@5 net@94 Clk net@78 Project1__nandBaseline
XnandBase@6 net@95 Clk net@79 Project1__nandBaseline
XnandBase@7 net@99 Clk net@80 Project1__nandBaseline
XnorBasel@0 net@37 net@0 net@4 Project1__norBaseline
XnorBasel@1 net@36 B net@4 Project1__norBaseline
XnorBasel@2 net@35 net@0 C Project1__norBaseline
XnorBasel@3 net@34 B C Project1__norBaseline
XnotBasel@0 B net@0 Project1__notBaseline
XnotBasel@1 C net@4 Project1__notBaseline
XnotBasel@2 net@73 net@77 Project1__notBaseline
XnotBasel@3 net@74 net@78 Project1__notBaseline
XnotBasel@5 net@76 net@80 Project1__notBaseline
Xwide_not@4 net@93 WL0 Project2__wide_not
Xwide_not@5 net@94 WL2 Project2__wide_not
Xwide_not@6 net@95 WL1 Project2__wide_not
Xwide_not@7 net@99 WL3 Project2__wide_not
.ENDS Project2__2_4_decoder

*** SUBCIRCUIT Project1__xorPass FROM CELL Project1:xorPass{sch}
.SUBCKT Project1__xorPass out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@150 y gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@166 net@130 net@150 gnd N L=0.022U W=0.022U
Mnmos@3 y x net@166 gnd N L=0.022U W=0.022U
Mnmos@4 net@130 x gnd gnd N L=0.022U W=0.022U
Mnmos@5 out net@166 gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd y net@150 vdd P L=0.022U W=0.022U
Mpmos@2 vdd x net@130 vdd P L=0.022U W=0.022U
Mpmos@3 vdd net@166 out vdd P L=0.022U W=0.022U
.ENDS Project1__xorPass

*** SUBCIRCUIT Project2__full_adder FROM CELL full_adder{sch}
.SUBCKT Project2__full_adder A B Cin Cout S
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@3 B A Project1__nandBaseline
XnandBase@1 net@16 net@17 Cin Project1__nandBaseline
XnandBase@2 Cout net@3 net@16 Project1__nandBaseline
XxorPass@0 net@17 B A Project1__xorPass
XxorPass@1 S Cin net@17 Project1__xorPass
.ENDS Project2__full_adder

*** SUBCIRCUIT Project2__deq_logic FROM CELL deq_logic{sch}
.SUBCKT Project2__deq_logic A A_next B B_next C C_next D
** GLOBAL gnd
** GLOBAL vdd
Xfull_add@0 C D gnd net@238 C_next Project2__full_adder
Xfull_add@1 B D net@238 net@243 B_next Project2__full_adder
Xfull_add@2 A D net@243 full_add@2_Cout A_next Project2__full_adder
.ENDS Project2__deq_logic

*** SUBCIRCUIT Project2__enq_logic FROM CELL enq_logic{sch}
.SUBCKT Project2__enq_logic A A_next B B_next C C_next E
** GLOBAL gnd
** GLOBAL vdd
Xfull_add@0 B E net@151 net@146 B_next Project2__full_adder
Xfull_add@1 C E gnd net@151 C_next Project2__full_adder
Xfull_add@2 A E net@146 full_add@2_Cout A_next Project2__full_adder
.ENDS Project2__enq_logic

*** SUBCIRCUIT Project2__and3 FROM CELL and3{sch}
.SUBCKT Project2__and3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@2 A net@11 gnd N L=0.022U W=0.022U
Mnmos@1 net@11 B net@12 gnd N L=0.022U W=0.022U
Mnmos@2 net@12 C gnd gnd N L=0.022U W=0.022U
Mnmos@3 O net@2 gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd C net@2 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@2 O vdd P L=0.022U W=0.022U
Mpmos@2 vdd B net@2 vdd P L=0.022U W=0.022U
Mpmos@3 vdd A net@2 vdd P L=0.022U W=0.022U
.ENDS Project2__and3

*** SUBCIRCUIT Project2__nor3 FROM CELL nor3{sch}
.SUBCKT Project2__nor3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O C gnd gnd N L=0.022U W=0.022U
Mnmos@1 O B gnd gnd N L=0.022U W=0.022U
Mnmos@2 O A gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A net@0 vdd P L=0.022U W=0.022U
Mpmos@1 net@0 B net@1 vdd P L=0.022U W=0.022U
Mpmos@2 net@1 C O vdd P L=0.022U W=0.022U
.ENDS Project2__nor3

*** SUBCIRCUIT Project2__size_logic FROM CELL size_logic{sch}
.SUBCKT Project2__size_logic A A_next B B_next C C_next D E Empty Full
** GLOBAL gnd
** GLOBAL vdd
Xand3@0 A B C Full Project2__and3
Xfull_add@0 C net@249 gnd net@158 C_next Project2__full_adder
Xfull_add@1 B net@245 net@158 net@163 B_next Project2__full_adder
Xfull_add@2 A net@245 net@163 full_add@2_Cout A_next Project2__full_adder
XnandBase@0 net@198 D net@199 Project1__nandBaseline
Xnor3@0 A B C Empty Project2__nor3
XnotBasel@3 net@198 net@245 Project1__notBaseline
XnotBasel@4 E net@199 Project1__notBaseline
XxorPass@0 net@249 D E Project1__xorPass
.ENDS Project2__size_logic

*** SUBCIRCUIT Project2__control_logic FROM CELL control_logic{sch}
.SUBCKT Project2__control_logic Clk D D_En DP_A DP_B DP_C E E_En Empty EP_A EP_B EP_C Full
** GLOBAL gnd
** GLOBAL vdd
Xdeq_logi@0 net@39 net@246 net@44 net@16 net@49 net@19 D_En Project2__deq_logic
Xenq_logi@0 net@54 net@257 net@59 net@9 net@64 net@12 E_En Project2__enq_logic
XnorBasel@0 D_En net@107 Empty Project1__norBaseline
XnorBasel@1 E_En net@106 Full Project1__norBaseline
XnotBasel@0 E net@106 Project1__notBaseline
XnotBasel@1 D net@107 Project1__notBaseline
XnotBasel@2 net@39 net@228 Project1__notBaseline
XnotBasel@3 net@44 net@232 Project1__notBaseline
XnotBasel@4 net@49 net@235 Project1__notBaseline
XnotBasel@5 net@54 net@240 Project1__notBaseline
XnotBasel@6 net@59 net@241 Project1__notBaseline
XnotBasel@7 net@64 net@242 Project1__notBaseline
Xregister@0 Clk net@246 net@39 HW7__register
Xregister@1 Clk net@16 net@44 HW7__register
Xregister@2 Clk net@19 net@49 HW7__register
Xregister@3 Clk net@257 net@54 HW7__register
Xregister@4 Clk net@9 net@59 HW7__register
Xregister@5 Clk net@12 net@64 HW7__register
Xregister@6 Clk net@266 net@69 HW7__register
Xregister@7 Clk net@2 net@74 HW7__register
Xregister@8 Clk net@5 net@79 HW7__register
Xsize_log@0 net@69 net@266 net@74 net@2 net@79 net@5 D_En E_En Empty Full Project2__size_logic
Xwide_not@1 net@228 DP_A Project2__wide_not
Xwide_not@6 net@232 DP_B Project2__wide_not
Xwide_not@7 net@235 DP_C Project2__wide_not
Xwide_not@8 net@240 EP_A Project2__wide_not
Xwide_not@9 net@241 EP_B Project2__wide_not
Xwide_not@10 net@242 EP_C Project2__wide_not
.ENDS Project2__control_logic

*** SUBCIRCUIT Project2__6TSRAM FROM CELL 6TSRAM{sch}
.SUBCKT Project2__6TSRAM BL BL_B R_WL W_WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Q W_WL BL gnd N L=0.022U W=0.22U
Mnmos@1 BL_B R_WL Qnot gnd N L=0.022U W=0.022U
Mnmos@2 Qnot Q gnd gnd N L=0.022U W=0.22U
Mnmos@3 Q Qnot gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd Q Qnot vdd P L=0.022U W=0.22U
Mpmos@1 vdd Qnot Q vdd P L=0.022U W=0.022U
.ENDS Project2__6TSRAM

*** SUBCIRCUIT Project2__word_cell FROM CELL word_cell{sch}
.SUBCKT Project2__word_cell BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL W_WL
** GLOBAL gnd
** GLOBAL vdd
X_6TSRAM@0 BL1_i BLB1_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@1 BL2_i BLB2_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@2 BL3_i BLB3_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@3 BL4_i BLB4_i R_WL W_WL Project2__6TSRAM
.ENDS Project2__word_cell

*** SUBCIRCUIT Project2__memory_block FROM CELL memory_block{sch}
.SUBCKT Project2__memory_block BL1_i BL2_i BL3_i BL4_i BL5_i BL6_i BL7_i BL8_i BLB1_i BLB2_i BLB3_i BLB4_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL1 R_WL2 R_WL3 R_WL4 W_WL1 W_WL2 W_WL3 W_WL4
** GLOBAL gnd
** GLOBAL vdd
Xword_cel@0 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL1 W_WL1 Project2__word_cell
Xword_cel@1 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL1 W_WL1 Project2__word_cell
Xword_cel@2 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL2 W_WL2 Project2__word_cell
Xword_cel@3 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL2 W_WL2 Project2__word_cell
Xword_cel@4 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL3 W_WL3 Project2__word_cell
Xword_cel@5 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL3 W_WL3 Project2__word_cell
Xword_cel@6 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL4 W_WL4 Project2__word_cell
Xword_cel@7 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL4 W_WL4 Project2__word_cell
.ENDS Project2__memory_block

*** SUBCIRCUIT Project2__precharge FROM CELL precharge{sch}
.SUBCKT Project2__precharge BL BL_B Clk_B
** GLOBAL vdd
Mpmos@0 vdd Clk_B BL_B vdd P L=0.022U W=0.022U
Mpmos@1 vdd Clk_B BL vdd P L=0.022U W=0.022U
.ENDS Project2__precharge

*** SUBCIRCUIT Project2__precharge_word FROM CELL precharge_word{sch}
.SUBCKT Project2__precharge_word BL1 BL2 BL3 BL4 BLB1 BLB2 BLB3 BLB4 Clk
** GLOBAL vdd
Xprecharg@0 BL1 BLB1 Clk Project2__precharge
Xprecharg@1 BL2 BLB2 Clk Project2__precharge
Xprecharg@2 BL3 BLB3 Clk Project2__precharge
Xprecharg@3 BL4 BLB4 Clk Project2__precharge
.ENDS Project2__precharge_word

*** SUBCIRCUIT Project2__tri_state_inverter FROM CELL tri_state_inverter{sch}
.SUBCKT Project2__tri_state_inverter data En Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@16 En gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@3 data gnd gnd N L=0.022U W=0.088U
Mnmos@2 net@3 En Out gnd N L=0.022U W=0.044U
Mpmos@0 vdd En net@16 vdd P L=0.022U W=0.022U
Mpmos@1 vdd data net@3 vdd P L=0.022U W=0.088U
Mpmos@2 Out net@16 net@3 vdd P L=0.022U W=0.044U
.ENDS Project2__tri_state_inverter

*** SUBCIRCUIT Project2__memory_core FROM CELL memory_core{sch}
.SUBCKT Project2__memory_core Clk_fast Clk_slow Deq Empty Enq Full I0 I1 I2 I3 O0 O1 O2 O3
** GLOBAL gnd
** GLOBAL vdd
X_2_4_deco@0 DB DC net@262 DEn net@16 net@17 net@18 net@19 Project2__2_4_decoder
X_2_4_deco@1 EB EC Clk_slow EEn net@20 net@21 net@22 net@23 Project2__2_4_decoder
Xcontrol_@0 Clk_slow Deq DEn DA DB DC Enq EEn Empty EA EB EC Full Project2__control_logic
Xmemory_b@0 WBL3 WBL2 WBL1 WBL0 WBL7 WBL6 WBL5 WBL4 RBL3 RBL2 RBL1 RBL0 RBL7 RBL6 RBL5 RBL4 net@16 net@17 net@18 net@19 net@20 net@21 net@22 net@23 Project2__memory_block
XnotBasel@0 EA net@66 Project1__notBaseline
XnotBasel@1 DA net@97 Project1__notBaseline
XnotBasel@2 Clk_slow net@262 Project1__notBaseline
Xprecharg@0 WBL3 WBL2 WBL1 WBL0 RBL3 RBL2 RBL1 RBL0 Clk_fast Project2__precharge_word
Xprecharg@1 WBL7 WBL6 WBL5 WBL4 RBL7 RBL6 RBL5 RBL4 Clk_fast Project2__precharge_word
Xtri_stat@1 I3 net@66 net@222 Project2__tri_state_inverter
Xtri_stat@2 I2 net@66 net@223 Project2__tri_state_inverter
Xtri_stat@3 I1 net@66 net@224 Project2__tri_state_inverter
Xtri_stat@4 I0 net@66 net@225 Project2__tri_state_inverter
Xtri_stat@5 I3 EA net@226 Project2__tri_state_inverter
Xtri_stat@6 I2 EA net@227 Project2__tri_state_inverter
Xtri_stat@7 I1 EA net@228 Project2__tri_state_inverter
Xtri_stat@8 I0 EA net@229 Project2__tri_state_inverter
Xtri_stat@9 RBL3 net@97 O3 Project2__tri_state_inverter
Xtri_stat@10 RBL2 net@97 O2 Project2__tri_state_inverter
Xtri_stat@11 RBL1 net@97 O1 Project2__tri_state_inverter
Xtri_stat@12 RBL0 net@97 O0 Project2__tri_state_inverter
Xtri_stat@13 RBL7 DA O3 Project2__tri_state_inverter
Xtri_stat@14 RBL6 DA O2 Project2__tri_state_inverter
Xtri_stat@15 RBL5 DA O1 Project2__tri_state_inverter
Xtri_stat@16 RBL4 DA O0 Project2__tri_state_inverter
Xvwide_no@0 net@222 WBL3 Project2__vwide_not
Xvwide_no@1 net@223 WBL2 Project2__vwide_not
Xvwide_no@2 net@224 WBL1 Project2__vwide_not
Xvwide_no@3 net@225 WBL0 Project2__vwide_not
Xvwide_no@4 net@226 WBL7 Project2__vwide_not
Xvwide_no@5 net@227 WBL6 Project2__vwide_not
Xvwide_no@6 net@228 WBL5 Project2__vwide_not
Xvwide_no@7 net@229 WBL4 Project2__vwide_not
.ENDS Project2__memory_core

.global gnd vdd

*** TOP LEVEL CELL: memory_core_test{sch}
VVPWL@0 Enq gnd pwl (0ns 0V .8ns 0V .9ns 1V 8.6ns 1V 8.7ns 0V) DC 0V AC 0V 0
VVPWL@1 Deq gnd pwl (0ns 0V 8.8ns 0V 8.9ns 1V 16.6ns 1V 16.7ns 0V) DC 0V AC 0V 0
VVPWL@2 I3 gnd pwl (0ns 0V 7.8ns 0V 7.9ns 1V 8.6ns 1V 8.7ns 0V) DC 0V AC 0V 0
VVPWL@3 I2 gnd pwl (0ns 0V 3.8ns 0V 3.9ns 1V 7.6ns 1V 7.7ns 0V) DC 0V AC 0V 0
VVPWL@4 I1 gnd pwl (0ns 0V 2.8ns 0V 2.9ns 1V 4.6ns 1V 4.7ns 0V 6.8ns 0V 6.9ns 1V 8.6ns 1V 8.7ns 0V) DC 0V AC 0V 0
VVPWL@5 I0 gnd pwl (0ns 0V .8ns 0V .9ns 1V 1.6ns 1V 1.7ns 0V 2.8ns 0V 2.9ns 1V 3.6ns 1V 3.7ns 0V 4.8ns 0V 4.9ns 1V 5.6ns 1V 5.7ns 0V 6.8ns 0V 6.9ns 1V 7.6ns 1V 7.7ns 0V) DC 0V AC 0V 0
VVPulse@0 Clk_double_freq gnd pulse (0 1V 0ns 0ps 0ps .5ns 1ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
Xclock_di@0 Clk_double_freq Clk Project2__clock_div
Xmemory_c@0 Clk_double_freq Clk Deq Empty Enq Full I0 I1 I2 I3 Out0 Out1 Out2 Out3 Project2__memory_core
.END
