*** SPICE deck for cell memory_core{sch} from library Project2
*** Created on Tue Dec 01, 2015 16:16:42
*** Last revised on Fri Dec 04, 2015 17:05:33
*** Written on Fri Dec 04, 2015 17:05:39 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /Users/neilnshah/Desktop/JUNIOR-YEAR/Fall15/Courses/ESE370/Project2/Project2/22nm_HP.pm

*** SUBCIRCUIT Project1__nandBaseline FROM CELL Project1:nandBaseline{sch}
.SUBCKT Project1__nandBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd x out vdd P L=0.022U W=0.022U
Mpmos@1 vdd y out vdd P L=0.022U W=0.022U
.ENDS Project1__nandBaseline

*** SUBCIRCUIT Project1__norBaseline FROM CELL Project1:norBaseline{sch}
.SUBCKT Project1__norBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x gnd gnd N L=0.022U W=0.022U
Mnmos@1 out y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd y net@10 vdd P L=0.022U W=0.022U
Mpmos@1 net@10 x out vdd P L=0.022U W=0.022U
.ENDS Project1__norBaseline

*** SUBCIRCUIT Project1__notBaseline FROM CELL Project1:notBaseline{sch}
.SUBCKT Project1__notBaseline in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd in out vdd P L=0.022U W=0.022U
.ENDS Project1__notBaseline

*** SUBCIRCUIT Project2__wide_not FROM CELL wide_not{sch}
.SUBCKT Project2__wide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.088U
Mpmos@0 vdd A O vdd P L=0.022U W=0.088U
.ENDS Project2__wide_not

*** SUBCIRCUIT Project2__2_4_decoder FROM CELL 2_4_decoder{sch}
.SUBCKT Project2__2_4_decoder B C En WL0 WL1 WL2 WL3
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@119 En net@37 Project1__nandBaseline
XnandBase@1 net@120 En net@36 Project1__nandBaseline
XnandBase@2 net@121 En net@35 Project1__nandBaseline
XnandBase@3 net@122 En net@34 Project1__nandBaseline
XnorBasel@0 net@37 B C Project1__norBaseline
XnorBasel@1 net@36 net@14 C Project1__norBaseline
XnorBasel@2 net@35 B net@23 Project1__norBaseline
XnorBasel@3 net@34 net@14 net@23 Project1__norBaseline
XnotBasel@2 C net@23 Project1__notBaseline
XnotBasel@3 B net@14 Project1__notBaseline
Xwide_not@4 net@119 WL0 Project2__wide_not
Xwide_not@5 net@120 WL2 Project2__wide_not
Xwide_not@6 net@121 WL1 Project2__wide_not
Xwide_not@7 net@122 WL3 Project2__wide_not
.ENDS Project2__2_4_decoder

*** SUBCIRCUIT Project1__xorPass FROM CELL Project1:xorPass{sch}
.SUBCKT Project1__xorPass out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 net@150 y gnd gnd N L=0.022U W=0.022U
Mnmos@2 net@166 net@130 net@150 gnd N L=0.022U W=0.022U
Mnmos@3 y x net@166 gnd N L=0.022U W=0.022U
Mnmos@4 net@130 x gnd gnd N L=0.022U W=0.022U
Mnmos@5 out net@166 gnd gnd N L=0.022U W=0.022U
Mpmos@1 vdd y net@150 vdd P L=0.022U W=0.022U
Mpmos@2 vdd x net@130 vdd P L=0.022U W=0.022U
Mpmos@3 vdd net@166 out vdd P L=0.022U W=0.022U
.ENDS Project1__xorPass

*** SUBCIRCUIT Project2__full_adder FROM CELL full_adder{sch}
.SUBCKT Project2__full_adder A B Cin Cout S
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@3 B A Project1__nandBaseline
XnandBase@1 net@16 net@17 Cin Project1__nandBaseline
XnandBase@2 Cout net@3 net@16 Project1__nandBaseline
XxorPass@0 net@17 B A Project1__xorPass
XxorPass@1 S Cin net@17 Project1__xorPass
.ENDS Project2__full_adder

*** SUBCIRCUIT Project2__deq_logic FROM CELL deq_logic{sch}
.SUBCKT Project2__deq_logic A A_next B B_next C C_next D
** GLOBAL gnd
** GLOBAL vdd
Xfull_add@0 C D gnd net@238 C_next Project2__full_adder
Xfull_add@1 B D net@238 net@243 B_next Project2__full_adder
Xfull_add@2 A D net@243 full_add@2_Cout A_next Project2__full_adder
.ENDS Project2__deq_logic

*** SUBCIRCUIT Project2__enq_logic FROM CELL enq_logic{sch}
.SUBCKT Project2__enq_logic A A_next B B_next C C_next E
** GLOBAL gnd
** GLOBAL vdd
Xfull_add@0 B E net@151 net@146 B_next Project2__full_adder
Xfull_add@1 C E gnd net@151 C_next Project2__full_adder
Xfull_add@2 A E net@146 full_add@2_Cout A_next Project2__full_adder
.ENDS Project2__enq_logic

*** SUBCIRCUIT HW7__nand_latch FROM CELL HW7:nand_latch{sch}
.SUBCKT HW7__nand_latch clock in out
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@0 in clock Project1__nandBaseline
XnandBase@1 net@11 a out Project1__nandBaseline
XnandBase@2 out net@0 net@11 Project1__nandBaseline
XnotBasel@0 clock a Project1__notBaseline
.ENDS HW7__nand_latch

*** SUBCIRCUIT HW7__register FROM CELL HW7:register{sch}
.SUBCKT HW7__register clock in out
** GLOBAL gnd
** GLOBAL vdd
Xnand_lat@0 clock mid out HW7__nand_latch
Xnand_lat@1 net@17 in mid HW7__nand_latch
XnotBasel@0 clock net@17 Project1__notBaseline
.ENDS HW7__register

*** SUBCIRCUIT Project2__and3 FROM CELL and3{sch}
.SUBCKT Project2__and3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@2 A net@11 gnd N L=0.022U W=0.022U
Mnmos@1 net@11 B net@12 gnd N L=0.022U W=0.022U
Mnmos@2 net@12 C gnd gnd N L=0.022U W=0.022U
Mnmos@3 O net@2 gnd gnd N L=0.022U W=0.088U
Mpmos@0 vdd C net@2 vdd P L=0.022U W=0.022U
Mpmos@1 vdd net@2 O vdd P L=0.022U W=0.088U
Mpmos@2 vdd B net@2 vdd P L=0.022U W=0.022U
Mpmos@3 vdd A net@2 vdd P L=0.022U W=0.022U
.ENDS Project2__and3

*** SUBCIRCUIT Project2__nor3 FROM CELL nor3{sch}
.SUBCKT Project2__nor3 A B C O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O C gnd gnd N L=0.022U W=0.022U
Mnmos@1 O B gnd gnd N L=0.022U W=0.022U
Mnmos@2 O A gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd A net@0 vdd P L=0.022U W=0.022U
Mpmos@1 net@0 B net@1 vdd P L=0.022U W=0.022U
Mpmos@2 net@1 C O vdd P L=0.022U W=0.022U
.ENDS Project2__nor3

*** SUBCIRCUIT Project2__nor4 FROM CELL nor4{sch}
.SUBCKT Project2__nor4 A B C D O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.022U
Mnmos@1 O B gnd gnd N L=0.022U W=0.022U
Mnmos@2 O C gnd gnd N L=0.022U W=0.022U
Mnmos@3 O D gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd D net@0 vdd P L=0.022U W=0.022U
Mpmos@1 net@0 C net@1 vdd P L=0.022U W=0.022U
Mpmos@2 net@1 B net@2 vdd P L=0.022U W=0.022U
Mpmos@3 net@2 A O vdd P L=0.022U W=0.022U
.ENDS Project2__nor4

*** SUBCIRCUIT Project2__size_logic FROM CELL size_logic{sch}
.SUBCKT Project2__size_logic D E Empty Full I0 I1 I2 I3 O0 O1 O2 O3
** GLOBAL gnd
** GLOBAL vdd
Xand3@1 net@265 net@266 net@269 net@245 Project2__and3
Xand3@2 net@269 net@296 net@266 net@250 Project2__and3
Xfull_add@0 I0 net@250 gnd net@158 O0 Project2__full_adder
Xfull_add@1 I1 net@245 net@158 net@163 O1 Project2__full_adder
Xfull_add@2 I2 net@245 net@163 net@301 O2 Project2__full_adder
Xfull_add@3 I3 net@245 net@301 full_add@3_Cout O3 Project2__full_adder
XnandBase@0 net@198 D net@199 Project1__nandBaseline
XnandBase@1 net@266 Full E Project1__nandBaseline
XnandBase@2 net@269 Empty D Project1__nandBaseline
XnandBase@4 net@321 net@348 I3 Project1__nandBaseline
Xnor3@0 I2 I1 I0 net@348 Project2__nor3
Xnor4@0 I2 I1 I0 I3 Empty Project2__nor4
XnotBasel@3 net@198 net@265 Project1__notBaseline
XnotBasel@4 E net@199 Project1__notBaseline
XnotBasel@5 net@321 Full Project1__notBaseline
XxorPass@0 net@296 D E Project1__xorPass
.ENDS Project2__size_logic

*** SUBCIRCUIT Project2__control_logic FROM CELL control_logic{sch}
.SUBCKT Project2__control_logic Clk D D_En DP_A DP_B DP_C E E_En Empty EP_A EP_B EP_C Full
** GLOBAL gnd
** GLOBAL vdd
Xdeq_logi@0 DPA net@246 DPB net@16 DPC net@19 D_En Project2__deq_logic
Xenq_logi@0 EPA net@257 EPB net@9 EPC net@12 E_En Project2__enq_logic
XnorBasel@0 D_En net@107 net@108 Project1__norBaseline
XnorBasel@1 E_En net@106 net@112 Project1__norBaseline
XnotBasel@0 E net@106 Project1__notBaseline
XnotBasel@1 D net@107 Project1__notBaseline
XnotBasel@2 DPA net@228 Project1__notBaseline
XnotBasel@3 DPB net@232 Project1__notBaseline
XnotBasel@4 DPC net@235 Project1__notBaseline
XnotBasel@5 EPA net@240 Project1__notBaseline
XnotBasel@6 EPB net@241 Project1__notBaseline
XnotBasel@7 EPC net@242 Project1__notBaseline
Xregister@0 Clk net@246 DPA HW7__register
Xregister@1 Clk net@16 DPB HW7__register
Xregister@2 Clk net@19 DPC HW7__register
Xregister@3 Clk net@257 EPA HW7__register
Xregister@4 Clk net@9 EPB HW7__register
Xregister@5 Clk net@12 EPC HW7__register
Xregister@6 Clk net@266 S3 HW7__register
Xregister@7 Clk net@2 S2 HW7__register
Xregister@8 Clk net@5 SC HW7__register
Xregister@9 Clk Full net@112 HW7__register
Xregister@10 Clk Empty net@108 HW7__register
Xregister@11 Clk net@291 S0 HW7__register
Xsize_log@0 D_En E_En Empty Full SC S2 S3 S0 net@5 net@2 net@266 net@291 Project2__size_logic
Xwide_not@1 net@228 DP_A Project2__wide_not
Xwide_not@6 net@232 DP_B Project2__wide_not
Xwide_not@7 net@235 DP_C Project2__wide_not
Xwide_not@8 net@240 EP_A Project2__wide_not
Xwide_not@9 net@241 EP_B Project2__wide_not
Xwide_not@10 net@242 EP_C Project2__wide_not
.ENDS Project2__control_logic

*** SUBCIRCUIT Project2__6TSRAM FROM CELL 6TSRAM{sch}
.SUBCKT Project2__6TSRAM BL BL_B R_WL W_WL
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 Q W_WL BL gnd N L=0.022U W=0.22U
Mnmos@1 BL_B R_WL Qnot gnd N L=0.022U W=0.022U
Mnmos@2 Qnot Q gnd gnd N L=0.022U W=0.22U
Mnmos@3 Q Qnot gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd Q Qnot vdd P L=0.022U W=0.22U
Mpmos@1 vdd Qnot Q vdd P L=0.022U W=0.022U
.ENDS Project2__6TSRAM

*** SUBCIRCUIT Project2__word_cell FROM CELL word_cell{sch}
.SUBCKT Project2__word_cell BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL W_WL
** GLOBAL gnd
** GLOBAL vdd
X_6TSRAM@0 BL1_i BLB1_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@1 BL2_i BLB2_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@2 BL3_i BLB3_i R_WL W_WL Project2__6TSRAM
X_6TSRAM@3 BL4_i BLB4_i R_WL W_WL Project2__6TSRAM
.ENDS Project2__word_cell

*** SUBCIRCUIT Project2__memory_block FROM CELL memory_block{sch}
.SUBCKT Project2__memory_block BL1_i BL2_i BL3_i BL4_i BL5_i BL6_i BL7_i BL8_i BLB1_i BLB2_i BLB3_i BLB4_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL1 R_WL2 R_WL3 R_WL4 W_WL1 W_WL2 W_WL3 W_WL4
** GLOBAL gnd
** GLOBAL vdd
Xword_cel@0 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL1 W_WL1 Project2__word_cell
Xword_cel@1 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL1 W_WL1 Project2__word_cell
Xword_cel@2 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL2 W_WL2 Project2__word_cell
Xword_cel@3 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL2 W_WL2 Project2__word_cell
Xword_cel@4 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL3 W_WL3 Project2__word_cell
Xword_cel@5 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL3 W_WL3 Project2__word_cell
Xword_cel@6 BL1_i BL2_i BL3_i BL4_i BLB1_i BLB2_i BLB3_i BLB4_i R_WL4 W_WL4 Project2__word_cell
Xword_cel@7 BL5_i BL6_i BL7_i BL8_i BLB5_i BLB6_i BLB7_i BLB8_i R_WL4 W_WL4 Project2__word_cell
.ENDS Project2__memory_block

*** SUBCIRCUIT Project2__precharge FROM CELL precharge{sch}
.SUBCKT Project2__precharge BL BL_B Clk_B
** GLOBAL vdd
Mpmos@0 vdd Clk_B BL_B vdd P L=0.022U W=0.44U
Mpmos@1 vdd Clk_B BL vdd P L=0.022U W=0.44U
.ENDS Project2__precharge

*** SUBCIRCUIT Project2__precharge_word FROM CELL precharge_word{sch}
.SUBCKT Project2__precharge_word BL1 BL2 BL3 BL4 BLB1 BLB2 BLB3 BLB4 Clk
** GLOBAL vdd
Xprecharg@0 BL1 BLB1 Clk Project2__precharge
Xprecharg@1 BL2 BLB2 Clk Project2__precharge
Xprecharg@2 BL3 BLB3 Clk Project2__precharge
Xprecharg@3 BL4 BLB4 Clk Project2__precharge
.ENDS Project2__precharge_word

*** SUBCIRCUIT Project2__tri_state_inverter FROM CELL tri_state_inverter{sch}
.SUBCKT Project2__tri_state_inverter data En Out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@16 En gnd gnd N L=0.022U W=0.022U
Mnmos@1 net@3 data gnd gnd N L=0.022U W=0.088U
Mnmos@2 net@3 En Out gnd N L=0.022U W=0.044U
Mpmos@0 vdd En net@16 vdd P L=0.022U W=0.022U
Mpmos@1 vdd data net@3 vdd P L=0.022U W=0.088U
Mpmos@2 Out net@16 net@3 vdd P L=0.022U W=0.044U
.ENDS Project2__tri_state_inverter

*** SUBCIRCUIT Project2__vvwide_not FROM CELL vvwide_not{sch}
.SUBCKT Project2__vvwide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.88U
Mpmos@0 vdd A O vdd P L=0.022U W=0.88U
.ENDS Project2__vvwide_not

*** SUBCIRCUIT Project2__vwide_not FROM CELL vwide_not{sch}
.SUBCKT Project2__vwide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.22U
Mpmos@0 vdd A O vdd P L=0.022U W=0.22U
.ENDS Project2__vwide_not

.global gnd vdd

*** TOP LEVEL CELL: memory_core{sch}
X_2_4_deco@0 DB DC DEn RWL0 RWL1 RWL2 RWL3 Project2__2_4_decoder
X_2_4_deco@1 EB EC EEn WWL0 WWL1 WWL2 wwl3_pre Project2__2_4_decoder
VVPWL@0 vpwl_wwl3 gnd pwl (0ns 0V 2.00ns 0V 2.01ns 1V 2.49ns 1V 2.50ns 0V 3.00ns 0V 3.01ns 1V 3.49ns 1V 3.50ns 0V) DC 0V AC 0V 0
Xcontrol_@0 Clk_slow Deq DEn DA DB DC Enq EEn Empty EA EB EC Full Project2__control_logic
Xmemory_b@0 WBL3 WBL2 WBL1 WBL0 WBL7 WBL6 WBL5 WBL4 RBL3 RBL2 RBL1 RBL0 RBL7 RBL6 RBL5 RBL4 RWL0 RWL1 RWL2 RWL3 WWL0 WWL1 WWL2 vpwl_wwl3 Project2__memory_block
XnandBase@0 wwl3_not wwl3_pre Clk_fast Project1__nandBaseline
XnotBasel@0 EA net@66 Project1__notBaseline
XnotBasel@1 DA net@97 Project1__notBaseline
XnotBasel@2 wwl3_not notBasel@2_out Project1__notBaseline
Xprecharg@0 WBL3 WBL2 WBL1 WBL0 RBL3 RBL2 RBL1 RBL0 Clk_fast Project2__precharge_word
Xprecharg@1 WBL7 WBL6 WBL5 WBL4 RBL7 RBL6 RBL5 RBL4 Clk_fast Project2__precharge_word
Xtri_stat@1 I3 net@66 net@280 Project2__tri_state_inverter
Xtri_stat@2 I2 net@66 net@281 Project2__tri_state_inverter
Xtri_stat@3 I1 net@66 net@282 Project2__tri_state_inverter
Xtri_stat@4 I0 net@66 net@283 Project2__tri_state_inverter
Xtri_stat@5 I3 EA net@284 Project2__tri_state_inverter
Xtri_stat@6 I2 EA net@285 Project2__tri_state_inverter
Xtri_stat@7 I1 EA net@286 Project2__tri_state_inverter
Xtri_stat@8 I0 EA net@287 Project2__tri_state_inverter
Xtri_stat@9 RBL3 net@97 O3 Project2__tri_state_inverter
Xtri_stat@10 RBL2 net@97 O2 Project2__tri_state_inverter
Xtri_stat@11 RBL1 net@97 O1 Project2__tri_state_inverter
Xtri_stat@12 RBL0 net@97 O0 Project2__tri_state_inverter
Xtri_stat@13 RBL7 DA O3 Project2__tri_state_inverter
Xtri_stat@14 RBL6 DA O2 Project2__tri_state_inverter
Xtri_stat@15 RBL5 DA O1 Project2__tri_state_inverter
Xtri_stat@16 RBL4 DA O0 Project2__tri_state_inverter
Xvvwide_n@0 net@295 WBL3 Project2__vvwide_not
Xvvwide_n@1 net@294 WBL2 Project2__vvwide_not
Xvvwide_n@2 net@293 WBL1 Project2__vvwide_not
Xvvwide_n@3 net@292 WBL0 Project2__vvwide_not
Xvvwide_n@4 net@291 WBL7 Project2__vvwide_not
Xvvwide_n@5 net@290 WBL6 Project2__vvwide_not
Xvvwide_n@6 net@289 WBL5 Project2__vvwide_not
Xvvwide_n@7 net@288 WBL4 Project2__vvwide_not
Xvwide_no@0 net@272 net@295 Project2__vwide_not
Xvwide_no@1 net@273 net@294 Project2__vwide_not
Xvwide_no@2 net@274 net@293 Project2__vwide_not
Xvwide_no@3 net@275 net@292 Project2__vwide_not
Xvwide_no@4 net@276 net@291 Project2__vwide_not
Xvwide_no@5 net@277 net@290 Project2__vwide_not
Xvwide_no@6 net@278 net@289 Project2__vwide_not
Xvwide_no@7 net@279 net@288 Project2__vwide_not
Xwide_not@16 net@280 net@272 Project2__wide_not
Xwide_not@17 net@281 net@273 Project2__wide_not
Xwide_not@18 net@282 net@274 Project2__wide_not
Xwide_not@19 net@283 net@275 Project2__wide_not
Xwide_not@20 net@284 net@276 Project2__wide_not
Xwide_not@21 net@285 net@277 Project2__wide_not
Xwide_not@22 net@286 net@278 Project2__wide_not
Xwide_not@23 net@287 net@279 Project2__wide_not
.END
