*** SPICE deck for cell 2_4_decoder_test{sch} from library Project2
*** Created on Thu Dec 03, 2015 22:52:37
*** Last revised on Thu Dec 03, 2015 22:58:47
*** Written on Thu Dec 03, 2015 23:05:25 by Electric VLSI Design System, version 9.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
* Model cards are described in this file:
.include /Users/neilnshah/Desktop/JUNIOR-YEAR/Fall15/Courses/ESE370/Project2/Project2/22nm_HP.pm

*** SUBCIRCUIT Project1__nandBaseline FROM CELL Project1:nandBaseline{sch}
.SUBCKT Project1__nandBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x net@13 gnd N L=0.022U W=0.022U
Mnmos@1 net@13 y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd x out vdd P L=0.022U W=0.022U
Mpmos@1 vdd y out vdd P L=0.022U W=0.022U
.ENDS Project1__nandBaseline

*** SUBCIRCUIT Project1__norBaseline FROM CELL Project1:norBaseline{sch}
.SUBCKT Project1__norBaseline out x y
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out x gnd gnd N L=0.022U W=0.022U
Mnmos@1 out y gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd y net@10 vdd P L=0.022U W=0.022U
Mpmos@1 net@10 x out vdd P L=0.022U W=0.022U
.ENDS Project1__norBaseline

*** SUBCIRCUIT Project1__notBaseline FROM CELL Project1:notBaseline{sch}
.SUBCKT Project1__notBaseline in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.022U W=0.022U
Mpmos@0 vdd in out vdd P L=0.022U W=0.022U
.ENDS Project1__notBaseline

*** SUBCIRCUIT Project2__wide_not FROM CELL wide_not{sch}
.SUBCKT Project2__wide_not A O
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 O A gnd gnd N L=0.022U W=0.088U
Mpmos@0 vdd A O vdd P L=0.022U W=0.088U
.ENDS Project2__wide_not

*** SUBCIRCUIT Project2__2_4_decoder FROM CELL 2_4_decoder{sch}
.SUBCKT Project2__2_4_decoder B C En WL0 WL1 WL2 WL3
** GLOBAL gnd
** GLOBAL vdd
XnandBase@0 net@119 En net@37 Project1__nandBaseline
XnandBase@1 net@120 En net@36 Project1__nandBaseline
XnandBase@2 net@121 En net@35 Project1__nandBaseline
XnandBase@3 net@122 En net@34 Project1__nandBaseline
XnorBasel@0 net@37 B C Project1__norBaseline
XnorBasel@1 net@36 net@14 C Project1__norBaseline
XnorBasel@2 net@35 B net@23 Project1__norBaseline
XnorBasel@3 net@34 net@14 net@23 Project1__norBaseline
XnotBasel@2 C net@23 Project1__notBaseline
XnotBasel@3 B net@14 Project1__notBaseline
Xwide_not@4 net@119 WL0 Project2__wide_not
Xwide_not@5 net@120 WL2 Project2__wide_not
Xwide_not@6 net@121 WL1 Project2__wide_not
Xwide_not@7 net@122 WL3 Project2__wide_not
.ENDS Project2__2_4_decoder

.global gnd vdd

*** TOP LEVEL CELL: 2_4_decoder_test{sch}
X_2_4_deco@0 B C En WL0 WL1 WL2 WL3 Project2__2_4_decoder
VVPulse@1 En gnd pulse (1V 0V 0ns 0ps 0ps 4ns 8ns) DC 0V AC 0V 0
VVPulse@2 C gnd pulse (1V 0V 0ns 0ps 0ps 1ns 2ns) DC 0V AC 0V 0
VVPulse@3 B gnd pulse (1V 0V 0ns 0ps 0ps 2ns 4ns) DC 0V AC 0V 0
VV_Generi@0 vdd gnd DC 1 AC 0
.END
